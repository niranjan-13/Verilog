`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:02:27 08/16/2022 
// Design Name: 
// Module Name:    dflipflop 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module dflipflop(
    input d,
    input clk,
    input rst,
    output reg q,
    output reg qb
    );
initial 
begin
q=1'b0;
qb=~q;
end
always@(posedge clk)
begin
if(rst)
q=0;
else
begin
case(d)
0:q=0;
1:q=1;
endcase
end
qb=~q;
end

endmodule
